---------------------------
--                       --
--         main          --
--                       --
---------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity main is
	port(
		BTN	:	in  std_logic_vector(0 downto 0);	-- Reset
		CLK	:	in  std_logic;				-- FPGA Clock
		
		-- Index sensor output
		LD	:	out std_logic_vector(1 downto 0);
		
		-- Index sensor
		JA2	:	in  std_logic;	-- Index 0
		JA8	:	in  std_logic;	-- Index 1
		
		-- Sensor 0
		JA9	:	in  std_logic;	-- HS1A		Motor 0 sensor 0
		JA3	:	in  std_logic;	-- HS1B		Motor 0 sensor 1
		
		-- Sensor 1
		JA4	:	in  std_logic;	-- HS2A		Motor 1 sensor 0
		JA10	:	in  std_logic;	-- HS2B		Motor 1 sensor 1
		
		-- Motor 0
		JB8	:	out std_logic;	-- ENA		Enable Motor 0
		JB3	:	out std_logic;	-- IN1A		Motor 0 pin 0
		JB9	:	out std_logic;	-- IN2A		Motor 0 pin 1
		
		-- Motor 1
		JB1	:	out std_logic;	-- ENA		Enable Motor 1
		JB2	:	out std_logic;	-- IN1B		Motor 1 pin 0
		JB7	:	out std_logic	-- IN2B		Motor 1 pin 1
		
		-- SPI0
		JC1	:	out std_logic;	-- SPI0CLK
		JC2	:	out std_logic;	-- SPI0SS
		JC3	:	out std_logic;	-- SPI0MOSI
		JC4	:	out std_logic;	-- SPI0MISO
		
		-- SPI1
		JC7	:	out std_logic;	-- SPI1CLK
		JC8	:	out std_logic;	-- SPI1SS
		JC9	:	out std_logic;	-- SPI1MOSI
		JC10	:	out std_logic	-- SPI1MISO
	);
end main;

architecture logic of main is
	
----------   Components   ----------
	
	component PWMController is
		generic(
			-- PWM Prescaler value
			constant PWMCLKScale	:	positive := 5;	-- Prescaled Clock = 50MHz / (PWMClockPrescaler * 2)
									-- PWMClockPrescaler -> 50MHz / (5 * 2) = 5MHz;
			-- PWM compare match bit width
			constant PWMBitWidth	:	positive := 8	-- PWM Frequency = 50MHz / (PWMClockPrescaler * 2 * (2 ** PWMBitWidth) - 4)
									-- PWM Frequency -> 50MHz / (5 * 2 * (2 ** 8) - 4) = 20KHz
		);
		port(
			RST		:	in  std_logic;
			CLK		:	in  std_logic;
		
			PWMCompareMatch	:	in  std_logic_vector((PWMBitWidth - 1) downto 0);
			PWMOutput	:	out std_logic_vector(1 downto 0)
		);
	end component;
	
begin
	
	-- Enable H-Bridge
	JB8 <= '1';
	
	PWMController0: PWMController
	generic map(
		PWMCLKScale => 5,	-- Prescaled Clock = 50MHz / (PWMClockPrescaler * 2)
					-- PWMClockPrescaler -> 50MHz / (5 * 2) = 5MHz;
		PWMBitWidth => 8	-- PWM Frequency = 50MHz / (PWMClockPrescaler * 2 * (2 ** PWMBitWidth) - 4)
					-- PWM Frequency -> 50MHz / (5 * 2 * (2 ** 8) - 4) = 20KHz
	)
	port map(
		RST => '0',
		CLK => CLK,
		PWMCompareMatch => SW(7 downto 0),
		PWMOutput(0) => JB3,
		PWMOutput(1) => JB9
	);
	
end logic;
